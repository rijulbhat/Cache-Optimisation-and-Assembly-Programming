library IEEE;
use IEEE.std_logic_1164.all;

entity test_decoder is
end entity;

architecture tb of test_decoder is
    signal alpha, beta, gamma, delta, en : std_logic;
    signal dec_output : std_logic_vector(15 downto 0);

    component decoder4x16 is 
    port(a, b, c, d, enable: in std_logic;
    dec: out std_logic_vector(15 downto 0));
    end component;

begin
    dut_instance: decoder4x16
    port map(a => alpha, b => beta, c => gamma, d => delta, enable => en, dec => dec_output);

    process 
    begin
        alpha <= '0';
        beta <= '0';
        gamma <= '0';
        delta <= '0';
        en <= '1';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '0';
        gamma <= '0';
        delta <= '1';
        en <= '1';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '0';
        gamma <= '1';
        delta <= '0';
        en <= '1';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '0';
        gamma <= '1';
        delta <= '1';
        en <= '1';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '1';
        gamma <= '0';
        delta <= '0';
        en <= '1';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '1';
        gamma <= '0';
        delta <= '1';
        en <= '1';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '1';
        gamma <= '1';
        delta <= '0';
        en <= '1';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '1';
        gamma <= '1';
        delta <= '1';
        en <= '1';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '0';
        gamma <= '0';
        delta <= '0';
        en <= '1';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '0';
        gamma <= '0';
        delta <= '1';
        en <= '1';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '0';
        gamma <= '1';
        delta <= '0';
        en <= '1';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '0';
        gamma <= '1';
        delta <= '1';
        en <= '1';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '1';
        gamma <= '0';
        delta <= '0';
        en <= '1';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '1';
        gamma <= '0';
        delta <= '1';
        en <= '1';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '1';
        gamma <= '1';
        delta <= '0';
        en <= '1';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '1';
        gamma <= '1';
        delta <= '1';
        en <= '1';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '0';
        gamma <= '0';
        delta <= '0';
        en <= '0';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '0';
        gamma <= '0';
        delta <= '1';
        en <= '0';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '0';
        gamma <= '1';
        delta <= '0';
        en <= '0';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '0';
        gamma <= '1';
        delta <= '1';
        en <= '0';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '1';
        gamma <= '0';
        delta <= '0';
        en <= '0';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '1';
        gamma <= '0';
        delta <= '1';
        en <= '0';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '1';
        gamma <= '1';
        delta <= '0';
        en <= '0';
        wait  for 1 ns;
        alpha <= '0';
        beta <= '1';
        gamma <= '1';
        delta <= '1';
        en <= '0';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '0';
        gamma <= '0';
        delta <= '0';
        en <= '0';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '0';
        gamma <= '0';
        delta <= '1';
        en <= '0';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '0';
        gamma <= '1';
        delta <= '0';
        en <= '0';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '0';
        gamma <= '1';
        delta <= '1';
        en <= '0';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '1';
        gamma <= '0';
        delta <= '0';
        en <= '0';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '1';
        gamma <= '0';
        delta <= '1';
        en <= '0';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '1';
        gamma <= '1';
        delta <= '0';
        en <= '0';
        wait  for 1 ns;
        alpha <= '1';
        beta <= '1';
        gamma <= '1';
        delta <= '1';
        en <= '0';
        wait  for 1 ns;
    end process;

end architecture;